module traffic_light_controller(red, yellow, red, car, clock, reset);
  input car
  input clock
  input reset
  output reg [1:0] red, yellow, green
 endmodule
